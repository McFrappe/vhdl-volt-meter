LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY lcd_full IS
	PORT
	(
		CLK :  IN  STD_LOGIC;
		RESET :  IN  STD_LOGIC;
		ENABLE :  IN  STD_LOGIC;
		DATA :  IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		LCD_RS :  OUT  STD_LOGIC;
		LCD_RW :  OUT  STD_LOGIC;
		LCD_ENABLE :  OUT  STD_LOGIC;
		LCD_BL :  OUT  STD_LOGIC;
		LCD_ON :  OUT  STD_LOGIC;
		LCD_BUSY :  OUT  STD_LOGIC;
		LCD_BUS :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END lcd_full;

ARCHITECTURE bdf_type OF lcd_full IS

COMPONENT lcd_controller
	PORT(CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 ENABLE : IN STD_LOGIC;
		 DATA : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 LCD_RS : OUT STD_LOGIC;
		 LCD_RW : OUT STD_LOGIC;
		 LCD_ENABLE : OUT STD_LOGIC;
		 LCD_BL : OUT STD_LOGIC;
		 LCD_ON : OUT STD_LOGIC;
		 LCD_BUSY : OUT STD_LOGIC;
		 LCD_BUS : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;



BEGIN



b2v_inst : lcd_controller
PORT MAP(CLK => CLK,
		 RESET => RESET,
		 ENABLE => ENABLE,
		 DATA => DATA,
		 LCD_RS => LCD_RS,
		 LCD_RW => LCD_RW,
		 LCD_ENABLE => LCD_ENABLE,
		 LCD_BL => LCD_BL,
		 LCD_ON => LCD_ON,
		 LCD_BUSY => LCD_BUSY,
		 LCD_BUS => LCD_BUS);


END bdf_type;